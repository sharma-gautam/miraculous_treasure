Miraculous Treasure
hello world
