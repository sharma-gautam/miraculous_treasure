Miraculous Treasure
